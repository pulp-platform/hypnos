//-----------------------------------------------------------------------------
// Title         : uCode Sequencer Package
//-----------------------------------------------------------------------------
// File          : pkg_ucode_sequencer.sv
// Author        : Manuel Eggimann  <meggimann@iis.ee.ethz.ch>
// Created       : 08.10.2018
//-----------------------------------------------------------------------------
// Description :
// Typedefinitions and parameters for the uCode Sequencer module.
//-----------------------------------------------------------------------------
// SPDX-License-Identifier: SHL-0.51
// Copyright (C) 2018-2021 ETH Zurich, University of Bologna
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License. You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//-----------------------------------------------------------------------------

package pkg_ucode_sequencer;
   import pkg_common::*;
   typedef logic [$clog2(ROWS_PER_HDVECT)-1:0] offset_t;

endpackage : pkg_ucode_sequencer
