//-----------------------------------------------------------------------------
// Title         : Definitions for module HD-Memory
//-----------------------------------------------------------------------------
// File          : pkg_hd_memory.sv
// Author        : Manuel Eggimann  <meggiman@blitzstein.ee.ethz.ch>
// Created       : 17.09.2018
//-----------------------------------------------------------------------------
// Description :
// 
//-----------------------------------------------------------------------------
// SPDX-License-Identifier: SHL-0.51 
// Copyright (C) 2018-2021 ETH Zurich, University of Bologna
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License. You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//-----------------------------------------------------------------------------

package pkg_hd_memory;
typedef   enum         logic[0:0] {WordMode, RowMode} write_mode_t;
endpackage : pkg_hd_memory
